module regfile(
    input         clk,
    // READ PORT 1
    input  [ 4:0] raddr1,
    output [31:0] rdata1,
    // READ PORT 2
    input  [ 4:0] raddr2,
    output [31:0] rdata2,
    // WRITE PORT
    input         rdt_req,
    input  [31:0] rdt_data,
    input  [ 4:0] rdt_addr,
    input         we,       //write enable, HIGH valid
    input  [ 4:0] waddr,
    input  [31:0] wdata
    `ifdef DIFFTEST_EN
    ,
    output [31:0] regs[31:0]
    `endif
);
reg [31:0] rf[31:0];
`ifdef DIFFTEST_EN
assign regs = rf;
`endif

//WRITE
always @(posedge clk) begin
    if (rdt_req) begin
        rf[rdt_addr] <= rdt_data;
        rf[waddr] <= wdata;
    end
    else if (we) rf[waddr]<= wdata;
end

//READ OUT 1
/* assign rdata1 = (raddr1==5'b0) ? 32'b0 : rf[raddr1]; */
assign rdata1 = {32{| raddr1}} & rf[raddr1]; //改动似乎不影响WNS

//READ OUT 2
/* assign rdata2 = (raddr2==5'b0) ? 32'b0 : rf[raddr2]; */
assign rdata2 = {32{| raddr2}} & rf[raddr2];

endmodule